module memory(
    input clk,
    input reset,
    input [7:0] data_in,
    output reg [7:0] data_out
);
   
	//место под запоминание
endmodule