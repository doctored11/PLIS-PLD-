module spiLedController(
    input clk,         
    input reset,        
    input inc,          
    input dec,          
    output SCLK,        
    output MOSI,        
    input MISO         
);
  
  //верхний уровень


endmodule