module counter(
    input clk,
    input reset,
    input inc,
    input dec,
    input [7:0] current_val,
    output reg [7:0] new_val
);
   //счетчик
endmodule