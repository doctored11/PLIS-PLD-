`timescale 1ns / 1ps
module spiLedController_tb();


endmodule