module spi_master(
    input clk,
    input [7:0] data,
    output reg SCLK,
    output reg MOSI,
    input MISO,
    output reg SS
);
   
	//реализация spi
endmodule