module spiLedController(
    input clk,         
    input reset,        
    input inc,          
    input dec,          
    output SCLK,        
    output MOSI,        
    input MISO         
);
  
  //верхний уровень
  /*
	 counter cnt(
			  .clk(clk),
			  .reset(reset),
			  .inc(inc),
			  .dec(dec),
			  .val(val)
		 );А
		 */

endmodule